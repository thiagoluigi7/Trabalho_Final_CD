module hexa7seg (digit0, digit1, LSD, MSD);
	input [3:0] digit0, digit1;
	output reg [6:0] LSD, MSD;
	
	always @*
	begin
		case(digit0)
			4'b0000: LSD <= 7'b0000001; // 0
			4'b0001: LSD <= 7'b1001111; // 1
			4'b0010: LSD <= 7'b0010010; // 2
			4'b0011: LSD <= 7'b0000110; // 3
			4'b0100: LSD <= 7'b1001100; // 4
			4'b0101: LSD <= 7'b0100100; // 5
			4'b0110: LSD <= 7'b0100000; // 6
			4'b0111: LSD <= 7'b0001111; // 7
			4'b1000: LSD <= 7'b0000000; // 8
			4'b1001: LSD <= 7'b0000100; // 9
			4'b1010: LSD <= 7'b0001000; // A
			4'b1011: LSD <= 7'b1100000; // b
			4'b1100: LSD <= 7'b0110001; // C
			4'b1101: LSD <= 7'b1000010; // d
			4'b1110: LSD <= 7'b0110000; // E
			4'b1111: LSD <= 7'b0111000; // F
		endcase 
			
		case(digit1)
			4'b0000: MSD <= 7'b0000001; // 0
			4'b0001: MSD <= 7'b1001111; // 1
			4'b0010: MSD <= 7'b0010010; // 2
			4'b0011: MSD <= 7'b0000110; // 3
			4'b0100: MSD <= 7'b1001100; // 4
			4'b0101: MSD <= 7'b0100100; // 5
			4'b0110: MSD <= 7'b0100000; // 6
			4'b0111: MSD <= 7'b0001111; // 7
			4'b1000: MSD <= 7'b0000000; // 8
			4'b1001: MSD <= 7'b0000100; // 9
			4'b1010: MSD <= 7'b0001000; // A
			4'b1011: MSD <= 7'b1100000; // b
			4'b1100: MSD <= 7'b0110001; // C
			4'b1101: MSD <= 7'b1000010; // d
			4'b1110: MSD <= 7'b0110000; // E
			4'b1111: MSD <= 7'b0111000; // F
		endcase
	
	end
	
endmodule
